*David Rubinstein
*class
*Assignment


*Netlist

*Sources

*Analysis


.op
.opt ingold=2 post

.end
